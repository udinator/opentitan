// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

class uart_sequencer extends dv_base_sequencer #(uart_item, uart_agent_cfg);
  `uvm_component_utils(uart_sequencer)

  `uvm_component_new

endclass
